// Карта памяти для модуля
localparam VERSION    = 32'h0000_0000; // RW
localparam DEBUG      = 32'h0000_0004; // RW
localparam FREQ_1     = 32'h0000_0008; // RW
localparam FREQ_2     = 32'h0000_000C; // RW
localparam FREQ_3     = 32'h0000_0010; // RW
localparam FREQ_4     = 32'h0000_0014; // RW
localparam FREQ_5     = 32'h0000_0018; // RW
localparam FREQ_6     = 32'h0000_001C; // RW
localparam FREQ_7     = 32'h0000_0020; // RW
localparam FREQ_8     = 32'h0000_0024; // RW
localparam FREQ_9     = 32'h0000_0028; // RW
localparam FREQ_10    = 32'h0000_002C; // RW
localparam FREQ_11    = 32'h0000_0030; // RW
localparam EN_CORDIC  = 32'h0000_0034; // RW
localparam STATUS     = 32'h0000_0038; // R 

